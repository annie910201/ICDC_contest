library verilog;
use verilog.vl_types.all;
entity CONV is
    generic(
        INITIAL         : integer := 0;
        READ_K0         : integer := 1;
        CONVOLUTION_K0  : integer := 2;
        RELU_K0         : integer := 3;
        WR_L0_K0        : integer := 4;
        RD_L0_K0        : integer := 5;
        WR_L1_K0        : integer := 6;
        READ_K1         : integer := 7;
        CONVOLUTION_K1  : integer := 8;
        RELU_K1         : integer := 9;
        WR_L0_K1        : integer := 10;
        RD_L0_K1        : integer := 11;
        WR_L1_K1        : integer := 12;
        BREAK_POINT     : integer := 13;
        RD_L1_K0        : integer := 14;
        WR_L2_K0        : integer := 15;
        RD_L1_K1        : integer := 16;
        WR_L2_K1        : integer := 17;
        FINISH          : integer := 18;
        K0_0            : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        K0_1            : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        K0_2            : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        K0_3            : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        K0_4            : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1);
        K0_5            : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        K0_6            : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        K0_7            : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        K0_8            : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        bias_0          : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        K1_0            : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        K1_1            : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        K1_2            : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        K1_3            : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1);
        K1_4            : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        K1_5            : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1);
        K1_6            : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        K1_7            : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1);
        K1_8            : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        bias_1          : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1)
    );
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        busy            : out    vl_logic;
        ready           : in     vl_logic;
        iaddr           : out    vl_logic_vector(11 downto 0);
        idata           : in     vl_logic_vector(19 downto 0);
        cwr             : out    vl_logic;
        caddr_wr        : out    vl_logic_vector(11 downto 0);
        cdata_wr        : out    vl_logic_vector(19 downto 0);
        crd             : out    vl_logic;
        caddr_rd        : out    vl_logic_vector(11 downto 0);
        cdata_rd        : in     vl_logic_vector(19 downto 0);
        csel            : out    vl_logic_vector(2 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of INITIAL : constant is 1;
    attribute mti_svvh_generic_type of READ_K0 : constant is 1;
    attribute mti_svvh_generic_type of CONVOLUTION_K0 : constant is 1;
    attribute mti_svvh_generic_type of RELU_K0 : constant is 1;
    attribute mti_svvh_generic_type of WR_L0_K0 : constant is 1;
    attribute mti_svvh_generic_type of RD_L0_K0 : constant is 1;
    attribute mti_svvh_generic_type of WR_L1_K0 : constant is 1;
    attribute mti_svvh_generic_type of READ_K1 : constant is 1;
    attribute mti_svvh_generic_type of CONVOLUTION_K1 : constant is 1;
    attribute mti_svvh_generic_type of RELU_K1 : constant is 1;
    attribute mti_svvh_generic_type of WR_L0_K1 : constant is 1;
    attribute mti_svvh_generic_type of RD_L0_K1 : constant is 1;
    attribute mti_svvh_generic_type of WR_L1_K1 : constant is 1;
    attribute mti_svvh_generic_type of BREAK_POINT : constant is 1;
    attribute mti_svvh_generic_type of RD_L1_K0 : constant is 1;
    attribute mti_svvh_generic_type of WR_L2_K0 : constant is 1;
    attribute mti_svvh_generic_type of RD_L1_K1 : constant is 1;
    attribute mti_svvh_generic_type of WR_L2_K1 : constant is 1;
    attribute mti_svvh_generic_type of FINISH : constant is 1;
    attribute mti_svvh_generic_type of K0_0 : constant is 1;
    attribute mti_svvh_generic_type of K0_1 : constant is 1;
    attribute mti_svvh_generic_type of K0_2 : constant is 1;
    attribute mti_svvh_generic_type of K0_3 : constant is 1;
    attribute mti_svvh_generic_type of K0_4 : constant is 1;
    attribute mti_svvh_generic_type of K0_5 : constant is 1;
    attribute mti_svvh_generic_type of K0_6 : constant is 1;
    attribute mti_svvh_generic_type of K0_7 : constant is 1;
    attribute mti_svvh_generic_type of K0_8 : constant is 1;
    attribute mti_svvh_generic_type of bias_0 : constant is 1;
    attribute mti_svvh_generic_type of K1_0 : constant is 1;
    attribute mti_svvh_generic_type of K1_1 : constant is 1;
    attribute mti_svvh_generic_type of K1_2 : constant is 1;
    attribute mti_svvh_generic_type of K1_3 : constant is 1;
    attribute mti_svvh_generic_type of K1_4 : constant is 1;
    attribute mti_svvh_generic_type of K1_5 : constant is 1;
    attribute mti_svvh_generic_type of K1_6 : constant is 1;
    attribute mti_svvh_generic_type of K1_7 : constant is 1;
    attribute mti_svvh_generic_type of K1_8 : constant is 1;
    attribute mti_svvh_generic_type of bias_1 : constant is 1;
end CONV;
